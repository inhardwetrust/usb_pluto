module ad936x_rx_to_axis(
    input [1:0] rx_data
    );
endmodule