module main(
    input  wire       clk,           // ????????? ????
    output reg  [0:0] interruptout,  // bit0 - ??? ?????
    output wire       inttest,        // ????? bit0 ?? ??????? ???
    output reg  [15:0] sample_out
);
    
    // --- ????????? ---
    // ??????? ?????? ??????? ?????????? reset ????? ??????:
    parameter integer POR_CYCLES     = 50_000_000;   // ~1 ??? ??? 50 ???
    // ?????? ????????: ?????? TOGGLE_CYCLES ?????? ?????? ??????? bit0
    parameter integer TOGGLE_CYCLES  = 10_000_000;   // ?? ????????? 1 ???

    // --- ?????????? reset (power-on) ---
    localparam integer POR_W = (POR_CYCLES > 1) ? $clog2(POR_CYCLES) : 1;
    reg [POR_W-1:0] por_cnt  = {POR_W{1'b0}};
    reg             rstn_loc = 1'b0;  // 0 ????? ????? ????????????

    always @(posedge clk) begin
        if (!rstn_loc) begin
            if (por_cnt == POR_CYCLES-1) begin
                rstn_loc <= 1'b1;               // ??????? reset
            end else begin
                por_cnt <= por_cnt + 1'b1;
            end
        end
    end

    // --- ???????? ??? ???????? bit0 ---
    localparam integer TG_W = (TOGGLE_CYCLES > 1) ? $clog2(TOGGLE_CYCLES) : 1;
    reg [TG_W-1:0] tg_cnt = {TG_W{1'b0}};
    reg            tog    = 1'b0;

    always @(posedge clk) begin
        if (!rstn_loc) begin
            tg_cnt       <= {TG_W{1'b0}};
            tog          <= 1'b0;
            interruptout <= 1'd0;
            
            sample_out<= 32'd866844501; ///sample_out<= 32'd866844501;
        end else begin
            if (tg_cnt == TOGGLE_CYCLES-1) begin
                tg_cnt <= {TG_W{1'b0}};
                tog    <= ~tog;                  // ????????? ?????? TOGGLE_CYCLES
            end else begin
                tg_cnt <= tg_cnt + 1'b1;
            end
            interruptout[0]   <= tog;
        end
    end

    assign inttest = interruptout[0];

endmodule
